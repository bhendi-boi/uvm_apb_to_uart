interface uart_intf ();
    logic rx_i;
    logic tx_o;
    logic event_o;
endinterface
