`define APB_ADDR_WIDTH 12
