`include "uvm_macros.svh"
`include "apb_intf.sv"

package apb_pkg;

    import uvm_pkg::*;
    `include "apb_types.sv"
    `include "apb_tr.sv"
    `include "apb_sequencer.sv"
    `include "apb_driver.sv"
    `include "apb_monitor.sv"
    `include "apb_coverage.sv"
    `include "apb_agent.sv"

    `include "apb_base_seq.sv"
    `include "apb_rand_seq.sv"

endpackage
